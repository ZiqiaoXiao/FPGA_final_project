module heart2_rom (
    input  wire        clk,
    input  wire [5:0]  pixel_x,
    input  wire [5:0]  pixel_y,
    output reg  [15:0] rgb_data
);
    reg [63:0] row_data;
    
   
    always @(*) begin
        case (pixel_y)
6'd0: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
 6'd1: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
 6'd2: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
 6'd3: row_data = 64'b0000011110011110000000000000000000000000000000000000000000000000;
 6'd4: row_data = 64'b0000111111111111100000000000000000000000000000000000000000000000;
 6'd5: row_data = 64'b0001111111111111111111111111111111111111111111111111111100000000;
 6'd6: row_data = 64'b0011111111111111111111111111111111111111111110000000000001100000;
 6'd7: row_data = 64'b0011111111111111111111111111111111111111111110000000000001100000;
 6'd8: row_data = 64'b0011111111111111111111111111111111111111111110000000000001100000;
 6'd9: row_data = 64'b0001111111111111111111111111111111111111111110000000000001100000;
6'd10: row_data = 64'b0000111111111111111111111111111111111111111110000000000001100000;
6'd11: row_data = 64'b0000011111111111111111111111111111111111111110000000000001100000;
6'd12: row_data = 64'b0000001111111111111111111111111111111111111111111111111110000000;
6'd13: row_data = 64'b0000000111111100000000000000000000000000000000000000000000000000;
6'd14: row_data = 64'b0000000011111000000000000000000000000000000000000000000000000000;
6'd15: row_data = 64'b0000000001100000000000000000000000000000000000000000000000000000;
6'd16: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd17: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd18: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd19: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;

        endcase
    end

    always @(posedge clk) begin
       
        rgb_data <= row_data[63-pixel_x] ? 16'hf800 : 16'h0000;
    end
endmodule