module start_rom (
    input  wire        clk,
    input  wire [5:0]  pixel_x,
    input  wire [5:0]  pixel_y,
    output reg  [15:0] rgb_data
);
    reg [63:0] row_data;
    
   
    always @(*) begin
        case (pixel_y)
6'd00: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd01: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd02: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd03: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd04: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd05: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd06: row_data = 64'b0000000000000000000000011111100000011111100000000000000000000000;
6'd07: row_data = 64'b0000000000000000000000100000011001100000010000000000000000000000;
6'd08: row_data = 64'b0000000000000000000001000000000110000000001000000000000000000000;
6'd09: row_data = 64'b0000000000000000000000100000001111000000010000000000000000000000;
6'd10: row_data = 64'b0000000000000000000000011011111001111101100000000000000000000000;
6'd11: row_data = 64'b0000000000000000000000000110001001000110000000000000000000000000;
6'd12: row_data = 64'b0000000000000000000000000000010000100000000000000000000000000000;
6'd13: row_data = 64'b0000000000000000000000000000010000100000000000000000000000000000;
6'd14: row_data = 64'b0000000000000000000000000000010000100000000000000000000000000000;
6'd15: row_data = 64'b0000000000000000000000000000110000110000000000000000000000000000;
6'd16: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd17: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd18: row_data = 64'b0000011111000111111111110000000100000001111111110001111111111100;
6'd19: row_data = 64'b0001110001100110011100110000000100000001111000111001100111001100;
6'd20: row_data = 64'b0011000000100100011100010000001110000001111000011101000111000100;
6'd21: row_data = 64'b0011100000000000011100000000001110000001111000011100000111000000;
6'd22: row_data = 64'b0011100000000000011100000000011011000001111000011100000111000000;
6'd23: row_data = 64'b0001111000000000011100000000011011000001111000011100000111000000;
6'd24: row_data = 64'b0001111110000000011100000000110001100001111000111000000111000000;
6'd25: row_data = 64'b0000111111100000011100000000110001100001111111100000000111000000;
6'd26: row_data = 64'b0000001111100000011100000001110001110001111011100000000111000000;
6'd27: row_data = 64'b0000000001110000011100000001111111110001111001110000000111000000;
6'd28: row_data = 64'b0000000000110000011100000011000000011001111001110000000111000000;
6'd29: row_data = 64'b0000000000110000011100000011000000011001111001111000000111000000;
6'd30: row_data = 64'b0011000000110000011100000011000000011001111000111000000111000000;
6'd31: row_data = 64'b0011100001100000011100000011000000011001111000111100000111000000;
6'd32: row_data = 64'b0000111111000000011100000111100000111101111000011100000111000000;
6'd33: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd34: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd35: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd36: row_data = 64'b0000000000000000000000000000011000000000000000000000000000000000;
6'd37: row_data = 64'b0000000000000000000000000001111111110000000000000000000000000000;
6'd38: row_data = 64'b0000000000000000110000000001100000111110000000000000000000000000;
6'd39: row_data = 64'b0000000000000000011111000000111000000111100000000000000000000000;
6'd40: row_data = 64'b0000000000000000000000111100000111000000111111000000000000000000;
6'd41: row_data = 64'b0000000000000000000000001111000001110000000111100000000000000000;
6'd42: row_data = 64'b0000000000000000000000000001111001100000000000000000000000000000;
6'd43: row_data = 64'b0000000000000000000000000000001111000000000000000000000000000000;
6'd44: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd45: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd46: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd47: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;



        endcase
    end

    always @(posedge clk) begin
        
        rgb_data <= row_data[63-pixel_x] ? 16'hFFE0 : 16'h0000;
    end
endmodule