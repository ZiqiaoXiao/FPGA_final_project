module win_rom (
    input  wire        clk,
    input  wire [5:0]  pixel_x,
    input  wire [5:0]  pixel_y,
    output reg  [15:0] rgb_data
);
    reg [63:0] row_data;
	 
	 
	 parameter C_BLACK  = 16'h0000;  
    parameter C_GREEN  = 16'h07E0;  
    parameter C_YELLOW = 16'hFFE0;  
    
    localparam Y_THRESHOLD = 6'd20;
    
    always @(*) begin
        case (pixel_y)
6'd00: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd01: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd02: row_data = 64'b0000011111000011111100001111100111110001111100000001111100000000;
6'd03: row_data = 64'b0000011111000011111100001111100111110001111110000001111100000000;
6'd04: row_data = 64'b0000011111000011111100001111100111110001111111000001111100000000;
6'd05: row_data = 64'b0000011111000011111100001111100111110001111101100001111100000000;
6'd06: row_data = 64'b0000011111000011111100001111100111110001111100110001111100000000;
6'd07: row_data = 64'b0000011111100011111100011111100111110001111100011001111100000000;
6'd08: row_data = 64'b0000001111110111111110111111000111110001111100001101111100000000;
6'd09: row_data = 64'b0000000111111110000111111110000111110001111100000111111100000000;
6'd10: row_data = 64'b0000000011111100000011111100000111110001111100000011111100000000;
6'd11: row_data = 64'b0000000011111100000011111100000111110001111100000001111100000000;
6'd12: row_data = 64'b0000000001111100000011111000000111110001111100000001111100000000;
6'd13: row_data = 64'b0000000001111100000011111000000111110001111100000001111100000000;
6'd14: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd15: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd16: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd17: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd18: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd19: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd20: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd21: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd22: row_data = 64'b0000000000000000000000000001111111111000000000000000000000000000;
6'd23: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
6'd24: row_data = 64'b0000000000000000000000000011111111111100000000000000000000000000;
6'd25: row_data = 64'b0000000000000000000000001101111111111011000000000000000000000000;
6'd26: row_data = 64'b0000000000000000000000010001111111111000100000000000000000000000;
6'd27: row_data = 64'b0000000000000000000000010001111111111000100000000000000000000000;
6'd28: row_data = 64'b0000000000000000000000001001111111111001000000000000000000000000;
6'd29: row_data = 64'b0000000000000000000000000111111111111110000000000000000000000000;
6'd30: row_data = 64'b0000000000000000000000000000011111110000000000000000000000000000;
6'd31: row_data = 64'b0000000000000000000000000000000110000000000000000000000000000000;
6'd32: row_data = 64'b0000000000000000000000000000000110000000000000000000000000000000;
6'd33: row_data = 64'b0000000000000000000000000000000110000000000000000000000000000000;
6'd34: row_data = 64'b0000000000000000000000000000011111100000000000000000000000000000;
6'd35: row_data = 64'b0000000000000000000000000111111111111110000000000000000000000000;
6'd36: row_data = 64'b0000000000000000000000000111111111111110000000000000000000000000;
6'd37: row_data = 64'b0000000000000000000000000111111111111110000000000000000000000000;
6'd38: row_data = 64'b0000000000000000000000000111111111111110000000000000000000000000;
6'd39: row_data = 64'b0000000000001111111111111111111111111110000000000000000000000000;
6'd40: row_data = 64'b0000000000001111111111111111111111111111111111111111110000000000;
6'd41: row_data = 64'b0000000000001111111111111111111111111111111111111111110000000000;
6'd42: row_data = 64'b0000000000001111111111111111111111111111111111111111110000000000;
6'd43: row_data = 64'b0000000000001111111111111111111111111111111111111111110000000000;
6'd44: row_data = 64'b0000000000001111111111111111111111111111111111111111110000000000;
6'd45: row_data = 64'b0000000000001111111111111111111111111111111111111111110000000000;
6'd46: row_data = 64'b0000000000001111111111111111111111111111111111111111110000000000;
6'd47: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;



        endcase
    end

    always @(posedge clk) begin
       
        if (row_data[63-pixel_x]) begin
            
            if (pixel_y <= Y_THRESHOLD) begin
                
                rgb_data <= C_GREEN; 
            end else begin
                
                rgb_data <= C_YELLOW; 
            end
        end else begin
           
            rgb_data <= C_BLACK;
        end
    end
endmodule