module emoji_rom (
    input  wire        clk,
    input  wire [5:0]  pixel_x,
    input  wire [5:0]  pixel_y,
    output reg  [15:0] rgb_data
);
    reg [63:0] row_data;
    
    parameter C_BLACK  = 16'h0000;
    parameter C_RED    = 16'hF800;
    parameter C_YELLOW = 16'hFFE0;
    
    localparam Y_START_RED = 6'd15;
    localparam Y_END_RED   = 6'd30;
    
    always @(*) begin
        case (pixel_y)
            6'd00: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd01: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd02: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd03: row_data = 64'b0000000000000000001111110000000001111110000000000000000000000000;
            6'd04: row_data = 64'b0000000000000000010000001110001110000001000000000000000000000000;
            6'd05: row_data = 64'b0000000000000000100000000001110000000000100000000000000000000000;
            6'd06: row_data = 64'b0000000000000000010000000011011000000001000000000000000000000000;
            6'd07: row_data = 64'b0000000000000000001111111010001011111110000000000000000000000000;
            6'd08: row_data = 64'b0000000000000000000000000110000100000000000000000000000000000000;
            6'd09: row_data = 64'b0000000000000000000000000110000110000000000000000000000000000000;
            6'd10: row_data = 64'b0000000000000000000000000110000110000000000000000000000000000000;
            6'd11: row_data = 64'b0000000000000000000000001100000110000000000000000000000000000000;
            6'd12: row_data = 64'b0000000000000000000000001000000001000000000000000000000000000000;
            6'd13: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd14: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd15: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd16: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd17: row_data = 64'b0000000011111111111100011100000000010001111111111100000000000000;
            6'd18: row_data = 64'b0000000011110000000000011110000000010001111000000011100000000000;
            6'd19: row_data = 64'b0000000011110000000000011111000000010001111000000001110000000000;
            6'd20: row_data = 64'b0000000011110000000000010111100000010001111000000001111000000000;
            6'd21: row_data = 64'b0000000011110000000000010011110000010001111000000000111100000000;
            6'd22: row_data = 64'b0000000011110000000000010001111000010001111000000000111100000000;
            6'd23: row_data = 64'b0000000011111111111100010000111100010001111000000000111100000000;
            6'd24: row_data = 64'b0000000011110000000000010000011110010001111000000000111100000000;
            6'd25: row_data = 64'b0000000011110000000000010000001111010001111000000000111100000000;
            6'd26: row_data = 64'b0000000011110000000000010000000111110001111000000001111100000000;
            6'd27: row_data = 64'b0000000011110000000000010000000011110001111000000001111000000000;
            6'd28: row_data = 64'b0000000011110000000000010000000001110001111000000011110000000000;
            6'd29: row_data = 64'b0000000011110000000000010000000000110001111000000111000000000000;
            6'd30: row_data = 64'b0000000011111111111100010000000000010001111111111000000000000000;
            6'd31: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd32: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd33: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd34: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd35: row_data = 64'b0000000000000000000000000000111110000000000000000000000000000000;
            6'd36: row_data = 64'b0000000000000000000000000011100011100000000000000000000000000000;
            6'd37: row_data = 64'b0000000000000111100000000111000001111110000000000000000000000000;
            6'd38: row_data = 64'b0000000000000001111110000011110000000111110000000000000000000000;
            6'd39: row_data = 64'b0000000000000000000111110000111111000000111111000000000000000000;
            6'd40: row_data = 64'b0000000000000000000000111111000001110000000011110000000000000000;
            6'd41: row_data = 64'b0000000000000000000000000011100011100000000000000000000000000000;
            6'd42: row_data = 64'b0000000000000000000000000000111110000000000000000000000000000000;
            6'd43: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd44: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd45: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd46: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd47: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd48: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd49: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd50: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd51: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd52: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd53: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd54: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd55: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd56: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd57: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd58: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd59: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd60: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd61: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd62: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
            6'd63: row_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        endcase
    end

    always @(posedge clk) begin
        if (row_data[63-pixel_x]) begin
            if (pixel_y >= Y_START_RED && pixel_y <= Y_END_RED) begin
                rgb_data <= C_RED; 
            end else begin
                rgb_data <= C_YELLOW; 
            end
        end else begin
            rgb_data <= C_BLACK;
        end
    end
endmodule